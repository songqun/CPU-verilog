`timescale 1ns / 1ps
module ssd(b, c);
	input [3:0] b;
	output reg [6:0] c;
	always @(b)
	begin
	case (b)
		4'b0000: c = ~7'b1111110;
		4'b0001: c = ~7'b0110000;
		4'b0010: c = ~7'b1101101;
		4'b0011: c = ~7'b1111001;
		4'b0100: c = ~7'b0110011;
		4'b0101: c = ~7'b1011011;
		4'b0110: c = ~7'b1011111;
		4'b0111: c = ~7'b1110000;
		4'b1000: c = ~7'b1111111;
		4'b1001: c = ~7'b1111011;
		4'b1010: c = ~7'b1110111;
		4'b1011: c = ~7'b0011111;
		4'b1100: c = ~7'b1001110;
		4'b1101: c = ~7'b0111101;
		4'b1110: c = ~7'b1001111;
		4'b1111: c = ~7'b1000111;
   endcase
	end
endmodule
